class trans;
  rand bit w_r;
  rand bit [7:0] data;
  rand bit [7:0] addr;
endclass
